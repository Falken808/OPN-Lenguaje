// Version del lenguaje OPN BluePanda

Version = 0.1.2
Release = V0.1.2
Name = OPN BluePanda
Codename = AutoVenv
Runtime = Python
CLI = opn
Features = venv_autogestion,pip_proxy,opn_json_dependencies,portable_build
